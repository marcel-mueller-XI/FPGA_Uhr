-- topClock fpga

