-- topClock

